//new project
